library ieee;
use ieee.std_logic_1164.all;

entity mux2x1_32Bits is
  -- Total de bits das entradas e saidas
  
  port (
    entradaA_MUX, entradaB_MUX   : in std_logic_vector(31 downto 0);
    seletor_MUX : in std_logic;
    saida_MUX : out std_logic_vector(31 downto 0)
  );
end entity;

architecture comportamento of mux2x1_32Bits is

  begin
  
    saida_MUX <= entradaA_MUX when (seletor_MUX = '0') else
					  entradaB_MUX when (seletor_MUX = '1');
					  
end architecture;