library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Baseado no apêndice C (Register Files) do COD (Patterson & Hennessy).

-- Entidade que define um banco de registradores com leitura de 2 registradores e escrita em 1 registrador simultaneamente.
entity bancoRegistradoresDiscretos is
    generic
    (
        larguraDados        : natural := 32;  -- Largura dos dados (em bits).
        larguraEndBancoRegs : natural := 5    -- Largura do endereço (2^5 = 32 posições).
    );
    port
    (
        clk        : in std_logic;  -- Sinal de clock.
        
        -- Entradas de endereços para os registradores de leitura (A e B) e de escrita (C).
        enderecoA  : in std_logic_vector((larguraEndBancoRegs-1) downto 0);
        enderecoB  : in std_logic_vector((larguraEndBancoRegs-1) downto 0);
        enderecoC  : in std_logic_vector((larguraEndBancoRegs-1) downto 0);

        -- Dado de escrita para o registrador C.
        dadoEscritaC : in std_logic_vector((larguraDados-1) downto 0);

        -- Sinal de controle de escrita. Se for '1', escreve no registrador C.
        escreveC  : in std_logic := '0';

        -- Saídas dos dados lidos dos registradores A e B.
        saidaA    : out std_logic_vector((larguraDados -1) downto 0);
        saidaB    : out std_logic_vector((larguraDados -1) downto 0)
    );
end entity bancoRegistradoresDiscretos;

-- Arquitetura comportamental do banco de registradores.
architecture comportamento of bancoRegistradoresDiscretos is

    -- Sinais auxiliares para lógica de bypass e seleção.
    signal bypassA, bypassB, zeroA, zeroB : std_logic;
    signal selectA, selectB : std_logic_vector(1 downto 0);
    
    -- Constante para representar o valor zero.
    constant zero : std_logic_vector(larguraDados-1 downto 0) := (others => '0');

    -- Sinais para armazenar os valores dos registradores.
    signal saidaReg0  : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg1  : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg2  : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg3  : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg4  : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg5  : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg6  : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg7  : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg8  : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg9  : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg10 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg11 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg12 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg13 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg14 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg15 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg16 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg17 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg18 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg19 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg20 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg21 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg22 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg23 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg24 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg25 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg26 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg27 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg28 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg29 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg30 : std_logic_vector(larguraDados-1 downto 0);
    signal saidaReg31 : std_logic_vector(larguraDados-1 downto 0);

    -- Sinais auxiliares para a lógica ENABLE de escrita.
    signal enableReg0  : std_logic;
    signal enableReg1  : std_logic;
    signal enableReg2  : std_logic;
    signal enableReg3  : std_logic;
    signal enableReg4  : std_logic;
    signal enableReg5  : std_logic;
    signal enableReg6  : std_logic;
    signal enableReg7  : std_logic;
    signal enableReg8  : std_logic;
    signal enableReg9  : std_logic;
    signal enableReg10 : std_logic;
    signal enableReg11 : std_logic;
    signal enableReg12 : std_logic;
    signal enableReg13 : std_logic;
    signal enableReg14 : std_logic;
    signal enableReg15 : std_logic;
    signal enableReg16 : std_logic;
    signal enableReg17 : std_logic;
    signal enableReg18 : std_logic;
    signal enableReg19 : std_logic;
    signal enableReg20 : std_logic;
    signal enableReg21 : std_logic;
    signal enableReg22 : std_logic;
    signal enableReg23 : std_logic;
    signal enableReg24 : std_logic;
    signal enableReg25 : std_logic;
    signal enableReg26 : std_logic;
    signal enableReg27 : std_logic;
    signal enableReg28 : std_logic;
    signal enableReg29 : std_logic;
    signal enableReg30 : std_logic;
    signal enableReg31 : std_logic;

    -- Saídas dos multiplexadores de seleção de registradores A e B.
    signal saida_mux32to1_A, saida_mux32to1_B : std_logic_vector(larguraDados-1 downto 0);
    
    -- Sinais para o resultado da operação XOR entre o endereço C e A/B.
    signal saida_muxEndC_XOR_EndA, saida_muxEndC_XOR_EndB : std_logic_vector(larguraDados-1 downto 0);
    
    -- Sinais para armazenar o resultado da operação XOR bit a bit entre C e A/B.
    signal xnorC_A : std_logic;
    signal xnorC_B : std_logic;

    -- Sinais para verificar se o endereço A ou B é zero.
    signal checa_Se_End_A_zero : std_logic;
    signal checa_Se_End_B_zero : std_logic;

begin

    -- Lógica para habilitar a escrita nos registradores baseados no endereço C.
    enableReg0  <= '1' when (escreveC = '1' and enderecoC = "00000") else '0';
    enableReg1  <= '1' when (escreveC = '1' and enderecoC = "00001") else '0';
    enableReg2  <= '1' when (escreveC = '1' and enderecoC = "00010") else '0';
    enableReg3  <= '1' when (escreveC = '1' and enderecoC = "00011") else '0';
    enableReg4  <= '1' when (escreveC = '1' and enderecoC = "00100") else '0';
    enableReg5  <= '1' when (escreveC = '1' and enderecoC = "00101") else '0';
    enableReg6  <= '1' when (escreveC = '1' and enderecoC = "00110") else '0';
    enableReg7  <= '1' when (escreveC = '1' and enderecoC = "00111") else '0';
    enableReg8  <= '1' when (escreveC = '1' and enderecoC = "01000") else '0';
    enableReg9  <= '1' when (escreveC = '1' and enderecoC = "01001") else '0';
    enableReg10 <= '1' when (escreveC = '1' and enderecoC = "01010") else '0';
    enableReg11 <= '1' when (escreveC = '1' and enderecoC = "01011") else '0';
    enableReg12 <= '1' when (escreveC = '1' and enderecoC = "01100") else '0';
    enableReg13 <= '1' when (escreveC = '1' and enderecoC = "01101") else '0';
    enableReg14 <= '1' when (escreveC = '1' and enderecoC = "01110") else '0';
    enableReg15 <= '1' when (escreveC = '1' and enderecoC = "01111") else '0';
    enableReg16 <= '1' when (escreveC = '1' and enderecoC = "10000") else '0';
    enableReg17 <= '1' when (escreveC = '1' and enderecoC = "10001") else '0';
    enableReg18 <= '1' when (escreveC = '1' and enderecoC = "10010") else '0';
    enableReg19 <= '1' when (escreveC = '1' and enderecoC = "10011") else '0';
    enableReg20 <= '1' when (escreveC = '1' and enderecoC = "10100") else '0';
    enableReg21 <= '1' when (escreveC = '1' and enderecoC = "10101") else '0';
    enableReg22 <= '1' when (escreveC = '1' and enderecoC = "10110") else '0';
    enableReg23 <= '1' when (escreveC = '1' and enderecoC = "10111") else '0';
    enableReg24 <= '1' when (escreveC = '1' and enderecoC = "11000") else '0';
    enableReg25 <= '1' when (escreveC = '1' and enderecoC = "11001") else '0';
    enableReg26 <= '1' when (escreveC = '1' and enderecoC = "11010") else '0';
    enableReg27 <= '1' when (escreveC = '1' and enderecoC = "11011") else '0';
    enableReg28 <= '1' when (escreveC = '1' and enderecoC = "11100") else '0';
    enableReg29 <= '1' when (escreveC = '1' and enderecoC = "11101") else '0';
    enableReg30 <= '1' when (escreveC = '1' and enderecoC = "11110") else '0';
    enableReg31 <= '1' when (escreveC = '1' and enderecoC = "11111") else '0';

    -- Instanciação dos 32 registradores genéricos (Reg0 até Reg31).
    Reg0 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg0, ENABLE => escreveC and enableReg0, CLK => clk, RST => '0');

    Reg1 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg1, ENABLE => escreveC and enableReg1, CLK => clk, RST => '0');

    Reg2 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg2, ENABLE => escreveC and enableReg2, CLK => clk, RST => '0');

    Reg3 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg3, ENABLE => escreveC and enableReg3, CLK => clk, RST => '0');

    Reg4 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg4, ENABLE => escreveC and enableReg4, CLK => clk, RST => '0');

    Reg5 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg5, ENABLE => escreveC and enableReg5, CLK => clk, RST => '0');

    Reg6 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg6, ENABLE => escreveC and enableReg6, CLK => clk, RST => '0');

    Reg7 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg7, ENABLE => escreveC and enableReg7, CLK => clk, RST => '0');

    Reg8 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg8, ENABLE => escreveC and enableReg8, CLK => clk, RST => '0');

    Reg9 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg9, ENABLE => escreveC and enableReg9, CLK => clk, RST => '0');

    Reg10 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg10, ENABLE => escreveC and enableReg10, CLK => clk, RST => '0');

    Reg11 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg11, ENABLE => escreveC and enableReg11, CLK => clk, RST => '0');

    Reg12 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg12, ENABLE => escreveC and enableReg12, CLK => clk, RST => '0');

    Reg13 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg13, ENABLE => escreveC and enableReg13, CLK => clk, RST => '0');

    Reg14 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg14, ENABLE => escreveC and enableReg14, CLK => clk, RST => '0');

    Reg15 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg15, ENABLE => escreveC and enableReg15, CLK => clk, RST => '0');

    Reg16 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg16, ENABLE => escreveC and enableReg16, CLK => clk, RST => '0');

    Reg17 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg17, ENABLE => escreveC and enableReg17, CLK => clk, RST => '0');

    Reg18 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg18, ENABLE => escreveC and enableReg18, CLK => clk, RST => '0');

    Reg19 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg19, ENABLE => escreveC and enableReg19, CLK => clk, RST => '0');

    Reg20 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg20, ENABLE => escreveC and enableReg20, CLK => clk, RST => '0');

    Reg21 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg21, ENABLE => escreveC and enableReg21, CLK => clk, RST => '0');

    Reg22 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg22, ENABLE => escreveC and enableReg22, CLK => clk, RST => '0');

    Reg23 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg23, ENABLE => escreveC and enableReg23, CLK => clk, RST => '0');

    Reg24 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg24, ENABLE => escreveC and enableReg24, CLK => clk, RST => '0');

    Reg25 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg25, ENABLE => escreveC and enableReg25, CLK => clk, RST => '0');

    Reg26 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg26, ENABLE => escreveC and enableReg26, CLK => clk, RST => '0');

    Reg27 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg27, ENABLE => escreveC and enableReg27, CLK => clk, RST => '0');

    Reg28 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg28, ENABLE => escreveC and enableReg28, CLK => clk, RST => '0');

    Reg29 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg29, ENABLE => escreveC and enableReg29, CLK => clk, RST => '0');

    Reg30 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg30, ENABLE => escreveC and enableReg30, CLK => clk, RST => '0');

    Reg31 : entity work.registradorGenerico
        generic map (larguraDados => larguraDados)
        port map (DIN => dadoEscritaC, DOUT => saidaReg31, ENABLE => escreveC and enableReg31, CLK => clk, RST => '0');

	 
	 mux32to1_A : entity work.mux32to1_32bits
		 generic map (LARGURA_DADOS => 32)
		 port map (
			  seletor => "00"& enderecoA,
			  saida => saida_mux32to1_A,
			  entrada0 => saidaReg0,
			  entrada1 => saidaReg1,
			  entrada2 => saidaReg2,
			  entrada3 => saidaReg3,
			  entrada4 => saidaReg4,
			  entrada5 => saidaReg5,
			  entrada6 => saidaReg6,
			  entrada7 => saidaReg7,
			  entrada8 => saidaReg8,
			  entrada9 => saidaReg9,
			  entrada10 => saidaReg10,
			  entrada11 => saidaReg11,
			  entrada12 => saidaReg12,
			  entrada13 => saidaReg13,
			  entrada14 => saidaReg14,
			  entrada15 => saidaReg15,
			  entrada16 => saidaReg16,
			  entrada17 => saidaReg17,
			  entrada18 => saidaReg18,
			  entrada19 => saidaReg19,
			  entrada20 => saidaReg20,
			  entrada21 => saidaReg21,
			  entrada22 => saidaReg22,
			  entrada23 => saidaReg23,
			  entrada24 => saidaReg24,
			  entrada25 => saidaReg25,
			  entrada26 => saidaReg26,
			  entrada27 => saidaReg27,
			  entrada28 => saidaReg28,
			  entrada29 => saidaReg29,
			  entrada30 => saidaReg30,
			  entrada31 => saidaReg31
		 );

	 xnorC_A <= '0' when 
		 ( enderecoA(0) XNOR enderecoC(0) ) AND
		 ( enderecoA(1) XNOR enderecoC(1) ) AND
		 ( enderecoA(2) XNOR enderecoC(2) ) --AND
		 --( enderecoA(3) XNOR enderecoC(3) ) AND
		 --( enderecoA(4) XNOR enderecoC(4) )
	else '1';
	
	 muxGenerico2x1_A : entity work.muxGenerico2x1
		 generic map (larguraDados => 32)
		 port map (
			  entradaA_MUX => dadoEscritaC,
			  entradaB_MUX => saida_mux32to1_A,
			  seletor_MUX => xnorC_A,
			  saida_MUX => saida_muxEndC_XOR_EndA
		 );
	
	checa_Se_End_A_zero <= '0' when (enderecoA = "00000") else '1';
	
	 mux_se_A_igual_0 : entity work.muxGenerico2x1
		 generic map (larguraDados => 32)
		 port map (
			  entradaA_MUX => x"00000000",
			  entradaB_MUX => saida_muxEndC_XOR_EndA,
			  seletor_MUX => checa_Se_End_A_zero,
			  saida_MUX => saidaA
		 );
	
	 mux32to1_B : entity work.mux32to1_32bits
		 generic map (LARGURA_DADOS => 32)
		 port map (
			  seletor => "00" & enderecoB,
			  saida => saida_mux32to1_B,
			  entrada0 => saidaReg0,
			  entrada1 => saidaReg1,
			  entrada2 => saidaReg2,
			  entrada3 => saidaReg3,
			  entrada4 => saidaReg4,
			  entrada5 => saidaReg5,
			  entrada6 => saidaReg6,
			  entrada7 => saidaReg7,
			  entrada8 => saidaReg8,
			  entrada9 => saidaReg9,
			  entrada10 => saidaReg10,
			  entrada11 => saidaReg11,
			  entrada12 => saidaReg12,
			  entrada13 => saidaReg13,
			  entrada14 => saidaReg14,
			  entrada15 => saidaReg15,
			  entrada16 => saidaReg16,
			  entrada17 => saidaReg17,
			  entrada18 => saidaReg18,
			  entrada19 => saidaReg19,
			  entrada20 => saidaReg20,
			  entrada21 => saidaReg21,
			  entrada22 => saidaReg22,
			  entrada23 => saidaReg23,
			  entrada24 => saidaReg24,
			  entrada25 => saidaReg25,
			  entrada26 => saidaReg26,
			  entrada27 => saidaReg27,
			  entrada28 => saidaReg28,
			  entrada29 => saidaReg29,
			  entrada30 => saidaReg30,
			  entrada31 => saidaReg31
		 );
	
	 xnorC_B <= '0' when 
		 ( enderecoB(0) XNOR enderecoC(0) ) AND
		 ( enderecoB(1) XNOR enderecoC(1) ) AND
		 ( enderecoB(2) XNOR enderecoC(2) ) --AND
		 --( enderecoB(3) XNOR enderecoC(3) ) AND
		 --( enderecoB(4) XNOR enderecoC(4) )
	else '1';
	
	 muxGenerico2x1_B : entity work.muxGenerico2x1
		 generic map (larguraDados => 32)
		 port map (
			  entradaA_MUX => dadoEscritaC,
			  entradaB_MUX => saida_mux32to1_B,
			  seletor_MUX => xnorC_B,
			  saida_MUX => saida_muxEndC_XOR_EndB
		 );
	
	 checa_Se_End_B_zero <= '0' when (enderecoB = "00000") else '1';
	
	 mux_se_B_igual_0 : entity work.muxGenerico2x1
		 generic map (larguraDados => 32)
		 port map (
			  entradaA_MUX => x"00000000",
			  entradaB_MUX => saida_muxEndC_XOR_EndB,
			  seletor_MUX => checa_Se_End_B_zero,
			  saida_MUX => saidaB
		 );

end architecture;
